* C:\Users\MohammadZakaria\Desktop\Semester-3rd-EEE\EEE-2302 Electronics Sessional\exp2\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Thu Feb 11 01:58:19 2021



** Analysis setup **
.tran 0ns 2ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
